@00000000
0010011100010000
1110110000010000
0000001000101011
1110001100001000
0111010100110000
1110110000010000
0000000000000100
1110001100001000
0000000000000000
1110110000010000
0000000000000001
1110001100001000
0100111000100000
1110110000010000
0000000000000010
1110001100001000
0000000000001010
1110110000010000
0000000000000011
1110001100001000
0000000000000001
1111110111001000
0000000000000010
1111110000010000
0000000000000011
1111010011010000
0000000000000010
1110001100001000
0000000000000010
1111110000010000
0000000000010100
1110001100000001
0110011111010001
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000000110
1110001100001000
0000011111010001
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000000111
1110001100001000
0111000011000001
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000001000101011
1111000010010000
0000000000001000
1110001100001000
0000011111010011
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000001001
1110001100001000
0110010001010010
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000001000101011
1111000010010000
0000000000001010
1110001100001000
0001010000110011
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000001011
1110001100001000
0110010100010110
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000001000101011
1111000010010000
0000000000001100
1110001100001000
0101101001101000
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000001101
1110001100001000
0110010100011010
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000001000101011
1111000010010000
0000000000001110
1110001100001000
0111110101000011
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000001000101011
1111000010010000
0000000000001111
1110001100001000
0111010100010010
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000001000101011
1111000010010000
0000000000010000
1110001100001000
0001100001100011
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000010001
1110001100001000
0110101101100010
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000010010
1110001100001000
0001011000110100
1110110000010000
0000000000000001
1111010011010000
0000000000000100
1111010011010000
0000000000010011
1110001100001000
0000000000000100
1111110010001000
1111110000010000
0000000000001000
1110001100000001
0100111000100000
1110110000010000
0000000000000000
1110001100001000